library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity single_cycle is
port(
    clk : in std_logic    
);
end entity single_cycle;

architecture structural of single_cycle is

begin

end architecture;
